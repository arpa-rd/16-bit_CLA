class transaction; 
  rand bit [15:0] a; 
  rand bit [15:0] b; 
  rand bit cin; 
  bit [15:0] sum; 
  bit cout; 
endclass:transaction 